// general_operation: General operation group
// Core Configuration Macros.
`define IOB_FUNCTIONS_VERSION 24'h008100
