// general_operation: General operation group
// Core Configuration Parameters Default Values
`define IOB_COUNTER_DATA_W 21
`define IOB_COUNTER_RST_VAL {DATA_W{1'b0}}
// Core Configuration Macros.
`define IOB_COUNTER_VERSION 24'h008100
