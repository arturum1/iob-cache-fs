// general_operation: General operation group
// Core Configuration Parameters Default Values
`define IOB_REG_CA_DATA_W 1
`define IOB_REG_CA_RST_VAL {DATA_W{1'b0}}
// Core Configuration Macros.
`define IOB_REG_CA_VERSION 24'h000100
