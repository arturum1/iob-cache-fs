// general_operation: General operation group
// Core Configuration Parameters Default Values
`define IOB_CACHE_CONTROL_DATA_W 32
`define IOB_CACHE_CONTROL_USE_CTRL_CNT 1
// Core Constants. DO NOT CHANGE
`define IOB_CACHE_CONTROL_VERSION 16'h0081
