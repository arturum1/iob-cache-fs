// general_operation: General operation group
// Core Configuration Parameters Default Values
`define IOB_RAM_T2P_HEXFILE "none"
`define IOB_RAM_T2P_ADDR_W 1
`define IOB_RAM_T2P_DATA_W 1
// Core Configuration Macros.
`define IOB_RAM_T2P_VERSION 24'h008100
