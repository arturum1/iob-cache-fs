// general_operation: General operation group
// Core Configuration Parameters Default Values
`define IOB_CACHE_IOB_CSRS_FE_ADDR_W 24
`define IOB_CACHE_IOB_CSRS_FE_DATA_W 32
`define IOB_CACHE_IOB_CSRS_BE_ADDR_W 24
`define IOB_CACHE_IOB_CSRS_BE_DATA_W 32
`define IOB_CACHE_IOB_CSRS_NWAYS_W 1
`define IOB_CACHE_IOB_CSRS_NLINES_W 7
`define IOB_CACHE_IOB_CSRS_WORD_OFFSET_W 3
`define IOB_CACHE_IOB_CSRS_WTBUF_DEPTH_W 4
`define IOB_CACHE_IOB_CSRS_REP_POLICY 0
`define IOB_CACHE_IOB_CSRS_WRITE_POL 0 
`define IOB_CACHE_IOB_CSRS_USE_CTRL 0
`define IOB_CACHE_IOB_CSRS_USE_CTRL_CNT 0
// Core Configuration Macros.
`define IOB_CACHE_IOB_CSRS_LRU 0
`define IOB_CACHE_IOB_CSRS_PLRU_MRU 1
`define IOB_CACHE_IOB_CSRS_PLRU_TREE 2
`define IOB_CACHE_IOB_CSRS_WRITE_THROUGH 0
`define IOB_CACHE_IOB_CSRS_WRITE_BACK 1
`define IOB_CACHE_IOB_CSRS_ADDR_W_CSRS 5
`define IOB_CACHE_IOB_CSRS_WTB_EMPTY_ADDR 0
`define IOB_CACHE_IOB_CSRS_WTB_EMPTY_W 8
`define IOB_CACHE_IOB_CSRS_WTB_FULL_ADDR 1
`define IOB_CACHE_IOB_CSRS_WTB_FULL_W 8
`define IOB_CACHE_IOB_CSRS_RW_HIT_ADDR 4
`define IOB_CACHE_IOB_CSRS_RW_HIT_W 32
`define IOB_CACHE_IOB_CSRS_RW_MISS_ADDR 8
`define IOB_CACHE_IOB_CSRS_RW_MISS_W 32
`define IOB_CACHE_IOB_CSRS_READ_HIT_ADDR 12
`define IOB_CACHE_IOB_CSRS_READ_HIT_W 32
`define IOB_CACHE_IOB_CSRS_READ_MISS_ADDR 16
`define IOB_CACHE_IOB_CSRS_READ_MISS_W 32
`define IOB_CACHE_IOB_CSRS_WRITE_HIT_ADDR 20
`define IOB_CACHE_IOB_CSRS_WRITE_HIT_W 32
`define IOB_CACHE_IOB_CSRS_WRITE_MISS_ADDR 24
`define IOB_CACHE_IOB_CSRS_WRITE_MISS_W 32
`define IOB_CACHE_IOB_CSRS_RST_CNTRS_ADDR 28
`define IOB_CACHE_IOB_CSRS_RST_CNTRS_W 8
`define IOB_CACHE_IOB_CSRS_INVALIDATE_ADDR 29
`define IOB_CACHE_IOB_CSRS_INVALIDATE_W 8
`define IOB_CACHE_IOB_CSRS_VERSION_ADDR 32
`define IOB_CACHE_IOB_CSRS_VERSION_W 32
`define IOB_CACHE_IOB_CSRS_VERSION 24'h000701
// Core Derived Parameters. DO NOT CHANGE
`define IOB_CACHE_IOB_CSRS_ADDR_W 6
`define IOB_CACHE_IOB_CSRS_FE_NBYTES FE_DATA_W / 8
`define IOB_CACHE_IOB_CSRS_FE_NBYTES_W $clog2(FE_NBYTES)
`define IOB_CACHE_IOB_CSRS_BE_NBYTES BE_DATA_W / 8
`define IOB_CACHE_IOB_CSRS_BE_NBYTES_W $clog2(BE_NBYTES)
`define IOB_CACHE_IOB_CSRS_LINE2BE_W WORD_OFFSET_W - $clog2(BE_DATA_W / FE_DATA_W)
`define IOB_CACHE_IOB_CSRS_DATA_W FE_DATA_W
