// general_operation: General operation group
// Core Configuration Parameters Default Values
`define IOB_CACHE_BACK_END_AXI_FE_ADDR_W 24
`define IOB_CACHE_BACK_END_AXI_FE_DATA_W 32
`define IOB_CACHE_BACK_END_AXI_BE_ADDR_W 24
`define IOB_CACHE_BACK_END_AXI_BE_DATA_W 32
`define IOB_CACHE_BACK_END_AXI_WORD_OFFSET_W 3
`define IOB_CACHE_BACK_END_AXI_WRITE_POL 0 
`define IOB_CACHE_BACK_END_AXI_AXI_ID_W 1
`define IOB_CACHE_BACK_END_AXI_AXI_ID 0
`define IOB_CACHE_BACK_END_AXI_AXI_LEN_W 4
`define IOB_CACHE_BACK_END_AXI_AXI_ADDR_W BE_ADDR_W
`define IOB_CACHE_BACK_END_AXI_AXI_DATA_W BE_DATA_W
// Core Configuration Macros.
`define IOB_CACHE_BACK_END_AXI_VERSION 24'h008100
// Core Derived Parameters. DO NOT CHANGE
`define IOB_CACHE_BACK_END_AXI_FE_NBYTES FE_DATA_W / 8
`define IOB_CACHE_BACK_END_AXI_FE_NBYTES_W $clog2(FE_NBYTES)
`define IOB_CACHE_BACK_END_AXI_BE_NBYTES BE_DATA_W / 8
`define IOB_CACHE_BACK_END_AXI_BE_NBYTES_W $clog2(BE_NBYTES)
`define IOB_CACHE_BACK_END_AXI_LINE2BE_W WORD_OFFSET_W - $clog2(BE_DATA_W / FE_DATA_W)
