// general_operation: General operation group
// Core Configuration Macros.
`define IOB_TASKS_VERSION 24'h008100
