// general_operation: General operation group
// Core Configuration Parameters Default Values
`define IOB_REGARRAY_SP_ADDR_W 2
`define IOB_REGARRAY_SP_DATA_W 21
// Core Constants. DO NOT CHANGE
`define IOB_REGARRAY_SP_VERSION 16'h0081
