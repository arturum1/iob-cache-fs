// general_operation: General operation group
// Core Configuration Parameters Default Values
`define IOB_RAM_SP_HEXFILE "none"
`define IOB_RAM_SP_DATA_W 8
`define IOB_RAM_SP_ADDR_W 14
// Core Configuration Macros.
`define IOB_RAM_SP_VERSION 24'h008100
// Core Derived Parameters. DO NOT CHANGE
`define IOB_RAM_SP_MEM_INIT_FILE_INT HEXFILE
