// general_operation: General operation group
// Core Constants. DO NOT CHANGE
`define IOB_TASKS_VERSION 16'h0081
