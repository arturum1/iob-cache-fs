//These macros may be dependent on instance parameters
//address macros
//addresses
`define IOB_CACHE_AXI_CSRS_WTB_EMPTY_ADDR 0
`define IOB_CACHE_AXI_CSRS_WTB_EMPTY_W 1

`define IOB_CACHE_AXI_CSRS_WTB_FULL_ADDR 1
`define IOB_CACHE_AXI_CSRS_WTB_FULL_W 1

`define IOB_CACHE_AXI_CSRS_RW_HIT_ADDR 4
`define IOB_CACHE_AXI_CSRS_RW_HIT_W 32

`define IOB_CACHE_AXI_CSRS_RW_MISS_ADDR 8
`define IOB_CACHE_AXI_CSRS_RW_MISS_W 32

`define IOB_CACHE_AXI_CSRS_READ_HIT_ADDR 12
`define IOB_CACHE_AXI_CSRS_READ_HIT_W 32

`define IOB_CACHE_AXI_CSRS_READ_MISS_ADDR 16
`define IOB_CACHE_AXI_CSRS_READ_MISS_W 32

`define IOB_CACHE_AXI_CSRS_WRITE_HIT_ADDR 20
`define IOB_CACHE_AXI_CSRS_WRITE_HIT_W 32

`define IOB_CACHE_AXI_CSRS_WRITE_MISS_ADDR 24
`define IOB_CACHE_AXI_CSRS_WRITE_MISS_W 32

`define IOB_CACHE_AXI_CSRS_RST_CNTRS_ADDR 28
`define IOB_CACHE_AXI_CSRS_RST_CNTRS_W 1

`define IOB_CACHE_AXI_CSRS_INVALIDATE_ADDR 29
`define IOB_CACHE_AXI_CSRS_INVALIDATE_W 1

`define IOB_CACHE_AXI_CSRS_VERSION_ADDR 30
`define IOB_CACHE_AXI_CSRS_VERSION_W 16

