// general_operation: General operation group
// Core Configuration Parameters Default Values
`define IOB_CACHE_IOB_CSRS_FE_ADDR_W 24
`define IOB_CACHE_IOB_CSRS_FE_DATA_W 32
`define IOB_CACHE_IOB_CSRS_BE_ADDR_W 24
`define IOB_CACHE_IOB_CSRS_BE_DATA_W 32
`define IOB_CACHE_IOB_CSRS_NWAYS_W 1
`define IOB_CACHE_IOB_CSRS_NLINES_W 7
`define IOB_CACHE_IOB_CSRS_WORD_OFFSET_W 3
`define IOB_CACHE_IOB_CSRS_WTBUF_DEPTH_W 4
`define IOB_CACHE_IOB_CSRS_REP_POLICY 0
`define IOB_CACHE_IOB_CSRS_WRITE_POL 0 
`define IOB_CACHE_IOB_CSRS_USE_CTRL 0
`define IOB_CACHE_IOB_CSRS_USE_CTRL_CNT 0
// Core Configuration Macros.
`define IOB_CACHE_IOB_CSRS_LRU 0
`define IOB_CACHE_IOB_CSRS_PLRU_MRU 1
`define IOB_CACHE_IOB_CSRS_PLRU_TREE 2
`define IOB_CACHE_IOB_CSRS_WRITE_THROUGH 0
`define IOB_CACHE_IOB_CSRS_WRITE_BACK 1
`define IOB_CACHE_IOB_CSRS_ADDR_W_CSRS 5
// Core Constants. DO NOT CHANGE
`define IOB_CACHE_IOB_CSRS_VERSION 16'h0071
// Core Derived Parameters. DO NOT CHANGE
`define IOB_CACHE_IOB_CSRS_ADDR_W 5
`define IOB_CACHE_IOB_CSRS_FE_NBYTES FE_DATA_W / 8
`define IOB_CACHE_IOB_CSRS_FE_NBYTES_W $clog2(FE_NBYTES)
`define IOB_CACHE_IOB_CSRS_BE_NBYTES BE_DATA_W / 8
`define IOB_CACHE_IOB_CSRS_BE_NBYTES_W $clog2(BE_NBYTES)
`define IOB_CACHE_IOB_CSRS_LINE2BE_W WORD_OFFSET_W - $clog2(BE_DATA_W / FE_DATA_W)
`define IOB_CACHE_IOB_CSRS_DATA_W FE_DATA_W
