// general_operation: General operation group
// Core Configuration Parameters Default Values
`define IOB_PRIO_ENC_W 21
`define IOB_PRIO_ENC_MODE "LOW"
// Core Configuration Macros.
`define IOB_PRIO_ENC_VERSION 24'h008100
