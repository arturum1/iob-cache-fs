// general_operation: General operation group
// Core Configuration Macros.
`define IOB_COVERAGE_ANALYZE_VERSION 24'h008100
